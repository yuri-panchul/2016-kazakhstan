module de0_cv
(
    input           CLOCK2_50,
    input           CLOCK3_50,
    inout           CLOCK4_50,
    input           CLOCK_50,
                   
    input           RESET_N,

    input   [ 3:0]  KEY,
    input   [ 9:0]  SW,

    output  [ 9:0]  LEDR,

    output  [ 6:0]  HEX0,
    output  [ 6:0]  HEX1,
    output  [ 6:0]  HEX2,
    output  [ 6:0]  HEX3,
    output  [ 6:0]  HEX4,
    output  [ 6:0]  HEX5,
                   
    output  [12:0]  DRAM_ADDR,
    output  [ 1:0]  DRAM_BA,
    output          DRAM_CAS_N,
    output          DRAM_CKE,
    output          DRAM_CLK,
    output          DRAM_CS_N,
    inout   [15:0]  DRAM_DQ,
    output          DRAM_LDQM,
    output          DRAM_RAS_N,
    output          DRAM_UDQM,
    output          DRAM_WE_N,
                   
    output  [ 3:0]  VGA_B,
    output  [ 3:0]  VGA_G,
    output          VGA_HS,
    output  [ 3:0]  VGA_R,
    output          VGA_VS,

    inout           PS2_CLK,
    inout           PS2_CLK2,
    inout           PS2_DAT,
    inout           PS2_DAT2,
                   
    output          SD_CLK,
    inout           SD_CMD,
    inout   [ 3:0]  SD_DATA,
                   
    inout   [35:0]  GPIO_0,
    inout   [35:0]  GPIO_1
);

    parameter [6:0] A = 7'b1110111,
                    L = 7'b1000111,
                    M = 7'b1101010,
                    N = 7'b0101010,
                    S = 7'b0010010,
                    T = 7'b0000111,
                    Y = 7'b0010001;

    wire sel = KEY [0];

    assign HEX5 =       A;
    assign HEX4 = sel ? L : S;
    assign HEX3 = sel ? M : T;
    assign HEX2 =       A;
    assign HEX1 = sel ? T : N;
    assign HEX0 = sel ? Y : A;

    // Alternative way
    
    // assign { HEX5, HEX4, HEX3, HEX2, HEX1, HEX0 } =
    //    sel ? { A, L, M, A, T, Y } : { A, S, T, A, N, A };

endmodule
